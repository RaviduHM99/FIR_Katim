package coeff_package is
    
end package coeff_package;